`ifndef _hhalfadder_h_
`define _hhalfadder_h_

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    03:47:40 08/07/2023 
// Design Name: 
// Module Name:    HalfAdder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module hHalfAdder(
    input a,
    input b,
	 output carry,
    output out
    );
	
	assign carry = a & b;
	assign out = a ^ b;

endmodule

`endif