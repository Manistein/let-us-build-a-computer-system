`ifndef _hub_v_ 
`define _hub_v_

module hub(
    input [15:0] instruction,
    input [15:0] pc_in,
    input is_loaded,

    output [15:0] pc_out
);



endmodule

`endif